NOM     | Prénom | Num. étudiant | Tél.              |  Mail                         |
--------------------------------------------------------------------------------------
JOFFRIN | Evan   | 22102052      | +33 6 07 68 15 07 |                               |
--------------------------------------------------------------------------------------
EL JAMAI| Ali    | 22104439      | +33 6 69 35 24 30 |                               |
--------------------------------------------------------------------------------------
PARIS   | Albin  | 22114221      |  06 14 90 74 81   |     paris.albin23@gmail.com   |
--------------------------------------------------------------------------------------
LEFORESTIER|Méril| 22104824      |  06 23 47 11 17   |meril.leforestier.3@gmail.com  |
--------------------------------------------------------------------------------------
BOURGUIBA |Adem        |22111078 |  07 81 14 79 38   | bourguibaaadem@yahoo.fr       |
--------------------------------------------------------------------------------------
ESPANET |   Nicolas | 22100628 |  06 49 40 12 29   | nicolas.espanet7@gmail.com      |
--------------------------------------------------------------------------------------
        |        |               |                   |                               |
--------------------------------------------------------------------------------------