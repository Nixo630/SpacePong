NOM     | Prénom | Num. étudiant | Tél.              |
------------------------------------------------------
JOFFRIN | Evan   | 22102052      | +33 6 07 68 15 07 |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------