NOM     | Prénom | Num. étudiant | Tél.              |
------------------------------------------------------
JOFFRIN | Evan   | 22102052      | +33 6 07 68 15 07 |
------------------------------------------------------
EL JAMAI| Ali    | 22104439      | +33 6 69 35 24 30 |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------
        |        |               |                   |
------------------------------------------------------