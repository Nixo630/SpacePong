NOM     | Prénom | Num. étudiant | Tél.              |  Mail                         |
--------------------------------------------------------------------------------------
JOFFRIN | Evan   | 22102052      | +33 6 07 68 15 07 |                               |
--------------------------------------------------------------------------------------
EL JAMAI| Ali    | 22104439      | +33 6 69 35 24 30 |                               |
--------------------------------------------------------------------------------------
PARIS   |Albin   | 22114221      |  06 14 90 74 81   |     paris.albin23@gmail.com   |
--------------------------------------------------------------------------------------
        |        |               |                   |                               |
--------------------------------------------------------------------------------------
        |        |               |                   |                               |
--------------------------------------------------------------------------------------
        |        |               |                   |                               |
--------------------------------------------------------------------------------------
        |        |               |                   |                               |
--------------------------------------------------------------------------------------